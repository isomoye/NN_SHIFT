module iverilog_dump();
initial begin
end
endmodule
